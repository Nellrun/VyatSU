-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II"
-- VERSION		"Version 9.1 Build 350 03/24/2010 Service Pack 2 SJ Web Edition"
-- CREATED		"Fri Oct 14 08:09:20 2011"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY aluip3 IS 
	PORT
	(
		S3 :  IN  STD_LOGIC;
		S2 :  IN  STD_LOGIC;
		M :  IN  STD_LOGIC;
		Cn :  IN  STD_LOGIC;
		S1 :  IN  STD_LOGIC;
		S0 :  IN  STD_LOGIC;
		A :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		B :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		Gn :  OUT  STD_LOGIC;
		Cn4 :  OUT  STD_LOGIC;
		Pn :  OUT  STD_LOGIC;
		AeqB :  OUT  STD_LOGIC;
		F :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END aluip3;

ARCHITECTURE bdf_type OF aluip3 IS 

SIGNAL	F_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_103 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_105 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_107 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_109 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_111 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;


BEGIN 
Gn <= SYNTHESIZED_WIRE_0;



SYNTHESIZED_WIRE_78 <= B(3) AND S3 AND A(3);


Cn4 <= NOT(SYNTHESIZED_WIRE_0 AND SYNTHESIZED_WIRE_1);


SYNTHESIZED_WIRE_5 <= SYNTHESIZED_WIRE_99 AND S1;


SYNTHESIZED_WIRE_6 <= S0 AND B(2);


SYNTHESIZED_WIRE_106 <= NOT(SYNTHESIZED_WIRE_3 OR SYNTHESIZED_WIRE_4);


SYNTHESIZED_WIRE_105 <= NOT(SYNTHESIZED_WIRE_5 OR SYNTHESIZED_WIRE_6 OR A(2));


SYNTHESIZED_WIRE_99 <= NOT(B(2));



SYNTHESIZED_WIRE_10 <= B(1) AND S3 AND A(1);


SYNTHESIZED_WIRE_9 <= A(1) AND S2 AND SYNTHESIZED_WIRE_100;


SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_100 AND S1;


SYNTHESIZED_WIRE_13 <= S0 AND B(1);


SYNTHESIZED_WIRE_108 <= NOT(SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10);


SYNTHESIZED_WIRE_77 <= A(3) AND S2 AND SYNTHESIZED_WIRE_101;


SYNTHESIZED_WIRE_107 <= NOT(SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13 OR A(1));


SYNTHESIZED_WIRE_100 <= NOT(B(1));



SYNTHESIZED_WIRE_17 <= B(0) AND S3 AND A(0);


SYNTHESIZED_WIRE_16 <= A(0) AND S2 AND SYNTHESIZED_WIRE_102;


SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_102 AND S1;


SYNTHESIZED_WIRE_19 <= S0 AND B(0);


SYNTHESIZED_WIRE_110 <= NOT(SYNTHESIZED_WIRE_16 OR SYNTHESIZED_WIRE_17);


SYNTHESIZED_WIRE_109 <= NOT(SYNTHESIZED_WIRE_18 OR SYNTHESIZED_WIRE_19 OR A(0));


SYNTHESIZED_WIRE_102 <= NOT(B(0));



SYNTHESIZED_WIRE_0 <= NOT(SYNTHESIZED_WIRE_103 OR SYNTHESIZED_WIRE_21 OR SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23);


SYNTHESIZED_WIRE_96 <= SYNTHESIZED_WIRE_101 AND S1;


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_104 AND SYNTHESIZED_WIRE_105;


SYNTHESIZED_WIRE_21 <= SYNTHESIZED_WIRE_104 AND SYNTHESIZED_WIRE_106 AND SYNTHESIZED_WIRE_107;


SYNTHESIZED_WIRE_23 <= SYNTHESIZED_WIRE_104 AND SYNTHESIZED_WIRE_106 AND SYNTHESIZED_WIRE_108 AND SYNTHESIZED_WIRE_109;


SYNTHESIZED_WIRE_1 <= NOT(SYNTHESIZED_WIRE_108 AND SYNTHESIZED_WIRE_106 AND SYNTHESIZED_WIRE_104 AND Cn AND SYNTHESIZED_WIRE_110 AND Cn);


Pn <= NOT(SYNTHESIZED_WIRE_104 AND SYNTHESIZED_WIRE_110 AND SYNTHESIZED_WIRE_106 AND SYNTHESIZED_WIRE_108);


SYNTHESIZED_WIRE_79 <= SYNTHESIZED_WIRE_108 AND Cn AND SYNTHESIZED_WIRE_110 AND SYNTHESIZED_WIRE_106 AND SYNTHESIZED_WIRE_111 AND SYNTHESIZED_WIRE_111;


SYNTHESIZED_WIRE_81 <= SYNTHESIZED_WIRE_108 AND SYNTHESIZED_WIRE_106 AND SYNTHESIZED_WIRE_109 AND SYNTHESIZED_WIRE_111;


SYNTHESIZED_WIRE_80 <= SYNTHESIZED_WIRE_106 AND SYNTHESIZED_WIRE_107 AND SYNTHESIZED_WIRE_111;


SYNTHESIZED_WIRE_82 <= SYNTHESIZED_WIRE_105 AND SYNTHESIZED_WIRE_111;


SYNTHESIZED_WIRE_85 <= Cn AND SYNTHESIZED_WIRE_110 AND SYNTHESIZED_WIRE_108 AND SYNTHESIZED_WIRE_111;


SYNTHESIZED_WIRE_97 <= S0 AND B(3);


SYNTHESIZED_WIRE_86 <= SYNTHESIZED_WIRE_108 AND SYNTHESIZED_WIRE_109 AND SYNTHESIZED_WIRE_111;


SYNTHESIZED_WIRE_87 <= SYNTHESIZED_WIRE_107 AND SYNTHESIZED_WIRE_111;


SYNTHESIZED_WIRE_93 <= Cn AND SYNTHESIZED_WIRE_110 AND SYNTHESIZED_WIRE_111;


SYNTHESIZED_WIRE_92 <= SYNTHESIZED_WIRE_109 AND SYNTHESIZED_WIRE_111;


SYNTHESIZED_WIRE_95 <= NOT(SYNTHESIZED_WIRE_111 AND Cn);


SYNTHESIZED_WIRE_83 <= SYNTHESIZED_WIRE_103 XOR SYNTHESIZED_WIRE_104;


SYNTHESIZED_WIRE_88 <= SYNTHESIZED_WIRE_106 XOR SYNTHESIZED_WIRE_105;


SYNTHESIZED_WIRE_90 <= SYNTHESIZED_WIRE_107 XOR SYNTHESIZED_WIRE_108;


SYNTHESIZED_WIRE_94 <= SYNTHESIZED_WIRE_109 XOR SYNTHESIZED_WIRE_110;


SYNTHESIZED_WIRE_111 <= NOT(M);



SYNTHESIZED_WIRE_104 <= NOT(SYNTHESIZED_WIRE_77 OR SYNTHESIZED_WIRE_78);


SYNTHESIZED_WIRE_84 <= NOT(SYNTHESIZED_WIRE_79 OR SYNTHESIZED_WIRE_80 OR SYNTHESIZED_WIRE_81 OR SYNTHESIZED_WIRE_82);


F_ALTERA_SYNTHESIZED(3) <= SYNTHESIZED_WIRE_83 XOR SYNTHESIZED_WIRE_84;


SYNTHESIZED_WIRE_89 <= NOT(SYNTHESIZED_WIRE_85 OR SYNTHESIZED_WIRE_86 OR SYNTHESIZED_WIRE_87);


F_ALTERA_SYNTHESIZED(2) <= SYNTHESIZED_WIRE_88 XOR SYNTHESIZED_WIRE_89;


F_ALTERA_SYNTHESIZED(1) <= SYNTHESIZED_WIRE_90 XOR SYNTHESIZED_WIRE_91;


SYNTHESIZED_WIRE_91 <= NOT(SYNTHESIZED_WIRE_92 OR SYNTHESIZED_WIRE_93);


F_ALTERA_SYNTHESIZED(0) <= SYNTHESIZED_WIRE_94 XOR SYNTHESIZED_WIRE_95;


AeqB <= F_ALTERA_SYNTHESIZED(0) AND F_ALTERA_SYNTHESIZED(1) AND F_ALTERA_SYNTHESIZED(2) AND F_ALTERA_SYNTHESIZED(3);


SYNTHESIZED_WIRE_103 <= NOT(SYNTHESIZED_WIRE_96 OR SYNTHESIZED_WIRE_97 OR A(3));


SYNTHESIZED_WIRE_101 <= NOT(B(3));



SYNTHESIZED_WIRE_4 <= B(2) AND S3 AND A(2);


SYNTHESIZED_WIRE_3 <= A(2) AND S2 AND SYNTHESIZED_WIRE_99;

F <= F_ALTERA_SYNTHESIZED;

END bdf_type;