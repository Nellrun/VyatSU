-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II"
-- VERSION		"Version 9.1 Build 350 03/24/2010 Service Pack 2 SJ Web Edition"
-- CREATED		"Thu Oct 13 14:47:38 2011"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY aluip4 IS 
	PORT
	(
		P4n :  IN  STD_LOGIC;
		P3n :  IN  STD_LOGIC;
		P2n :  IN  STD_LOGIC;
		P1n :  IN  STD_LOGIC;
		G4n :  IN  STD_LOGIC;
		G3n :  IN  STD_LOGIC;
		G2n :  IN  STD_LOGIC;
		G1n :  IN  STD_LOGIC;
		Cn :  IN  STD_LOGIC;
		Pn :  OUT  STD_LOGIC;
		Gn :  OUT  STD_LOGIC;
		Cz :  OUT  STD_LOGIC;
		Cy :  OUT  STD_LOGIC;
		Cx :  OUT  STD_LOGIC
	);
END aluip4;

ARCHITECTURE bdf_type OF aluip4 IS 

SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;


BEGIN 



Pn <= NOT(SYNTHESIZED_WIRE_39 AND SYNTHESIZED_WIRE_40 AND SYNTHESIZED_WIRE_41 AND SYNTHESIZED_WIRE_42);


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_39 AND SYNTHESIZED_WIRE_41 AND SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_43;


Gn <= NOT(SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10 OR SYNTHESIZED_WIRE_11);


Cz <= SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13 OR SYNTHESIZED_WIRE_44 OR SYNTHESIZED_WIRE_15;


Cy <= SYNTHESIZED_WIRE_16 OR SYNTHESIZED_WIRE_45 OR SYNTHESIZED_WIRE_18;


Cx <= SYNTHESIZED_WIRE_43 OR SYNTHESIZED_WIRE_20;


SYNTHESIZED_WIRE_39 <= NOT(P4n);



SYNTHESIZED_WIRE_41 <= NOT(P3n);



SYNTHESIZED_WIRE_42 <= NOT(P2n);



SYNTHESIZED_WIRE_40 <= NOT(P1n);



SYNTHESIZED_WIRE_11 <= NOT(G4n);



SYNTHESIZED_WIRE_10 <= SYNTHESIZED_WIRE_39 AND SYNTHESIZED_WIRE_41 AND SYNTHESIZED_WIRE_45;


SYNTHESIZED_WIRE_44 <= NOT(G3n);



SYNTHESIZED_WIRE_45 <= NOT(G2n);



SYNTHESIZED_WIRE_43 <= NOT(G1n);



SYNTHESIZED_WIRE_9 <= SYNTHESIZED_WIRE_39 AND SYNTHESIZED_WIRE_44;


SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_41 AND SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_40 AND Cn;


SYNTHESIZED_WIRE_15 <= SYNTHESIZED_WIRE_41 AND SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_43;


SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_41 AND SYNTHESIZED_WIRE_45;


SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_40 AND Cn;


SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_43;


SYNTHESIZED_WIRE_20 <= SYNTHESIZED_WIRE_40 AND Cn;


END bdf_type;