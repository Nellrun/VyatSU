library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_encoder is

	port
	(
		addr	: in natural range 0 to 256;
		clk		: in std_logic;
		q		: out std_logic_vector(3 downto 0)
	);
	
end entity;

architecture rtl of rom_encoder is

	-- Build a 2-D array type for the RoM
	subtype word_t is std_logic_vector(3 downto 0);
	type memory_t is array(255 downto 0) of word_t;
		
	function init_rom
		return memory_t is
		variable tmp : memory_t := (others => (others => '0'));
		begin
			for addr_pos in 0 to 256 loop
				-- Initialize each address with the address itself
				tmp(addr_pos) := std_logic_vector(to_unsigned(addr_pos, 4));
			end loop;
		return tmp;
	end init_rom;
	
	-- Declare the ROM signal and specify a default value.	Quartus II
	-- will create a memory initialization file (.mif) based on the 
	-- default value.
	signal rom : memory_t := (
		0 => "0000",
		1 => "0001",
		2 => "0010",
		4 => "0011",
		8 => "0100",
		16 => "0101",
		32 => "0110",
		64 => "0111",
		128 => "1000",
		OTHERS => "0000"
	);
	
begin
	
	process(clk)
	begin
		if(rising_edge(clk)) then
			q <= rom(addr);
		end if;
	end process;
		
end rtl;
